* ADA4530 Macro-model
* Function: Operational Amplifier
*
* Revision History:
* Rev 0 Oct 2015: ZF/VW
* Tested by PN at Vsy=+/-5V
* Copyright 2015 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spicemodels/license
* for License Statement. Use of this model indicates your acceptance
* of the terms and provisions in the License Staement.
*
* Guard output pins GRD1, GRD2 should be left unconnected for simulation purpose.
* DNC pin should be left unconnected for simulation purpose.
* Tested on MultSIm, SiMetrix(NGSpice), PSpice.
*
* Not modeled: Distortion, PSRR, Overload Recovery,
*              Shutdown Turn On/Turn Off time.
*
* Parameters (typical values) modeled include:
*   Vos, Ibias, Input CM limits and Typ output voltge swing,
*   Open Loop Gain & Phase, Slew Rate, Output current limits, Voltage & Current Noise,
*   Capacitive load drive, supply currents, supply functionality.
*
* Not simulated/implemented - performance over temp
* Parameter variations with supply are not modeled
*
* CAUTION!!  
* To aid in convergence, most Spice simulators add a
* conductance on every node to insure that no node is floating.
* This is GMIN, and the default value is usually 1E-12.  To properly 
* simulate the low input bias current and low current noise, the 
* Spice simulator options have to be set to the following:
* GMIN=1E-16
* ABSTOL=1E-16
* RSHUNT=1E16 (Multisim)
*
* When using model in Multisim, comment out the first .ends ADA4530 statement
* and uncomment the second .ends ADA4530 statement.
*
* In some simulations, number of iterations (ITL1) may have to be increased to aid convergence.
*
*
*
* Node Assignments
*                Non-Inverting Input
*                |   Inverting Input
*                |    |    Positive supply
*                |    |    |    Negative supply
*                |    |    |    |    Output
*                |    |    |    |    |    GRD1
*                |    |    |    |    |    |    GRD2
*                |    |    |    |    |    |    |
*.Subckt ADA4530 N100 N101 N102 N103 N104 N105 N106
.Subckt ADA4530_3rdparty_ver N100 N101 N102 N103 N104 N105 N106
*
X1	N100	N101	N102	N103	1	Amplifier
X2	N100	2	N102	N103	3	Buffer
R1	1	N104	Rideal	20
R2	2	3	Rideal	1e-6
R3	3	4	Rideal	1e3
R4	4	N105	Rideal	1e-6
R5	4	N106	Rideal	1e-6
R6	N105	0	Rideal	1e9
R7	N106	0	Rideal	1e9
.model	Rideal	res(T_ABS=-273)
*
* .ends ada4530 
*
*
**********************************************
.Subckt Amplifier 100 101 102 103 104
**********************************************
***Power Supplies***
Rz	102	1020	Rideal	10
DzPS	98	1020	diode
S1	98	103	106	113	Switch
R1	1020	99	Rideal	1e7
R2	99	103	Rideal	1e7
e1	111	110	1020	110	1
e2	110	112	110	103	1
e3	110	0	99	0	1
*
*
***Inputs***
VOS	100	2	dc	8e-6
IbiasP	110	2	dc	1e-15
IbiasN	110	101	dc	1e-15
*RinCMP	110	2	Rideal	100e12
*RinCMN	9	110	Rideal	100e12
CinCMP	110	2	2.4e-12
CinCMN	101	110	2.4e-12
IOS	101	2	1e-15
*RinDiff	9	2	Rideal	100e12
CinDiff	101	2	0.6e-12
EVN 9 0 101 0 1
*
*
***Non-Inverting Input with Clamp***
g1	3	110	110	2	0.001
RInP	3	110	Rideal	1e3
RX1	40	3	Rideal	1
DInP	40	41	diode
DInN	42	40	diode
VinP	111	41	dc	1.96
VinN	42	112	dc	0.46
*
*
***Vnoise***
hVn	6	5	Vmeas1	707.10678
Vmeas1	20	110	DC	0
Vvn	21	110	dc	0.65
Dvn	21	20	DVnoisy
hVn1	6	7	Vmeas2	707.10678
Vmeas2	22	110	dc	0
Vvn1	23	110	dc	0.65
Dvn1	23	22	DVnoisy
*
*
***Inoise***
FnIN	9	110	Vmeas3	0.7071068
Vmeas3	51	110	dc	0
VnIN	50	110	dc	0.65
DnIN	50	51	DINnoisy
FnIN1	110	9	Vmeas4	0.7071068
Vmeas4	53	110	dc	0
VnIN1	52	110	dc	0.65
DnIN1	52	53	DINnoisy
*
FnIP	2	110	Vmeas5	0.7071068
Vmeas5	31	110	dc	0
VnIP	30	110	dc	0.65
DnIP	30	31	DIPnoisy
FnIP1	110	2	Vmeas6	0.7071068
Vmeas6	33	110	dc	0
VnIP1	32	110	dc	0.65
DnIP1	32	33	DIPnoisy
*
*
***CMRR***
RcmrrP	3	10	Rideal	1e12
RcmrrN	10	9	Rideal	1e12
g10	11	110	10	110	-9e-8
Lcmrr	11	12	1e-12
Rcmrr	12	110	Rideal	1e3
e4	5	3	11	110	1
*
*
***Power Down***
VPD	111	80	dc	0.8
VPD1	81	0	dc	0.1
RPD	111	106	Rideal	1e6
ePD	80	113	82	0	1
RDP1	82	0	Rideal	1e3
CPD	82	0	1e-10
S5	81	82	83	113	Switch
CDP1	83	0	1e-12
RPD2	106	83	1e6
*
*
***Gain Split***
g200	200	110	7	9	1
R200	200	110	Rideal	1e5
*
*
***Dominant Pole at 0.14 Hz***
g210	210	110	Value={limit(V(200,110)*1.242e-5,.1413,-.1413)}
R210	210	110	Rideal	1.137e7
C210	210	110	1e-7
*
*
***Output Voltage Clamp-1***
RX2	60	210	Rideal	0.001
DzVoutP	61	60	DzVoutP
DzVoutN	60	62	DzVoutN
DVoutP	61	63	diode
DVoutN	64	62	diode
VoutP	65	63	dc	5.03
VoutN	64	66	dc	5.015
e60	65	110	111	110	1.014
e61	66	110	112	110	1.114
*
*
***Pole at 17MHz***
g220	220	110	210	110	0.001
R220	220	110	Rideal	1000
C220	220	110	9.362e-12
*
***Pole at 40MHz***
g230	230	110	220	110	0.001
R230	230	110	Rideal	1000
C230	230	110	3.9789e-12
*
***Pole at 40MHz***
g240	240	110	230	110	0.001
R240	240	110	Rideal	1000
C240	240	110	3.9789e-12
*
***Pole at 45MHz***
g245	245	110	240	110	0.001
R245	245	110	Rideal	1000
C245	245	110	3.5368e-12
*
***Pole at 45MHz***
g250	250	110	245	110	0.001
R250	250	110	Rideal	1000
C250	250	110	3.5368e-12
*
***Pole at 45MHz***
g255	255	110	250	110	0.001
R255	255	110	Rideal	1000
C255	255	110	3.5368e-12
*
***Pole at 50MHz***
g260	260	110	255	110	0.001
R260	260	110	Rideal	1000
C260	260	110	3.1831e-12
*
***Pole at 50MHz***
g265	265	110	260	110	0.001
R265	265	110	Rideal	1000
C265	265	110	3.1831e-12
*
***Pole at 50MHz***
g270	270	110	265	110	0.001
R270	270	110	Rideal	1000
C270	270	110	3.1831e-12
*
***Notch: f=12MHz, Zeta=0.7, Gain=2.5dB***
e280	280	110	270	110	1
L280	285	281	378.78e-9
C280	281	282	464.398e-12
R281	282	110	Rideal	29.983
R280	280	285	Rideal	10
*
***Peak: f=9MHz, Zeta=1, Gain=2.7dB***
e290	290	110	285	110	1
L290	290	291	88.419e-9
C290	291	292	3536.773e-12
R291	292	110	Rideal	27.429
e295	295	110	292	110	1.3646
R290	290	292	Rideal	10
*
*
***Output Stage***
g300	300	110	295	110	0.001
R300	300	110	Rideal	1000
e301	301	110	300	110	1
Rout	302	303	Rideal	 90
Lout	303	310	 3700e-9
Cout	310	110	 16e-12
*
*
***Output Current Limit***
H1	301	304	Vsense1	100
Vsense1	301	302	dc	0
VIoutP	305	304	dc	0.836
VIoutN	304	306	dc	2.336
DIoutP	307	305	diode
DIoutN	306	307	diode
Rx3	307	300	Rideal	100
*
*
***Output Clamp-2***
VoutP1	111	73	dc	0.7
VoutN1	74	112	dc	0.7102
DVoutP1	75	73	diode
DVoutN1	74	75	diode
RX4	75	310	Rideal	0.001
*
*
***Supply Currents***
FIoVcc	314	110	Vmeas8	1
Vmeas8	310	311	dc	0
R314	110	314	Rideal	1e9
DzOVcc	110	314	diode
DOVcc	102	314	diode
RX5	311	312	Rideal	0.001
FIoVee	315	110	Vmeas9	1
Vmeas9	312	313	dc	0
R315	315	110	Rideal	1e9
DzOVee	315	110	diode
DOVee	315	103	diode
*
*
***Output Switch***
S4	104	313	106	113	Switch
*
*
*** Common Models ***
.model	diode	d(bv=100)
.model	Switch	vswitch(Von=0.15,Voff=0.05,ron=10,roff=1e6)
.model	DzVoutP	D(BV=4.3)
.model	DzVoutN	D(BV=4.3)
.model	DzSlewP	D(BV=13.546)
.model	DzSlewN	D(BV=13.546)
.model	DVnoisy	D(IS=7.28e-15 KF=8.83e-17)
.model	DINnoisy	D(IS=1.87e-25 KF=0)
.model	DIPnoisy	D(IS=1.87e-25 KF=0)
.model	Rideal	res(T_ABS=-273)
*
.ends Amplifier
*
*
**********************************************
.Subckt Buffer 100 101 102 103 104
**********************************************
***Power Supplies***
Rz1	102	1020	Rideal	10
Rz2	103	1030	Rideal	10
R3	96	0	Rideal	1e3
S6	97	96	1020	1030	Sswitch
V2	97	0	dc	2
gBias	1020	1030	96	0	0.09e-3
DzPS	98	1020	diode
gQuies	1020	98	96	0	0.81e-3
S1	98	1030	106	113	Switch
R1	1020	99	Rideal	1e7
R2	99	1030	Rideal	1e7
e1	111	110	1020	110	1
e2	110	112	110	1030	1
e3	110	0	99	0	1
*
*
***Inputs***
S2	1	100	106	113	Switch
S3	9	101	106	113	Switch
VOS	1	2	dc	0
*IbiasP	110	2	dc	0
*IbiasN	110	9	dc	0
*RinCMP	110	2	Rideal	100e12
*RinCMN	9	110	Rideal	100e12
CinCMP	110	2	1e-15
CinCMN	9	110	1e-15
*IOS	9	2	0
*RinDiff	9	2	Rideal	100e12
CinDiff	9	2	1e-15
*
*
***Non-Inverting Input with Clamp***
g1	3	110	110	2	0.001
RInP	3	110	Rideal	1e3
RX1	40	3	Rideal	1
DInP	40	41	diode
DInN	42	40	diode
VinP	111	41	dc	1.96
VinN	42	112	dc	0.56
*
*
***Vnoise***
hVn	6	5	Vmeas1	707.10678
Vmeas1	20	110	DC	0
Vvn	21	110	dc	0.65
Dvn	21	20	DVnoisy
hVn1	6	7	Vmeas2	707.10678
Vmeas2	22	110	dc	0
Vvn1	23	110	dc	0.65
Dvn1	23	22	DVnoisy
*
*
***Inoise***
FnIN	9	110	Vmeas3	0.7071068
Vmeas3	51	110	dc	0
VnIN	50	110	dc	0.65
DnIN	50	51	DINnoisy
FnIN1	110	9	Vmeas4	0.7071068
Vmeas4	53	110	dc	0
VnIN1	52	110	dc	0.65
DnIN1	52	53	DINnoisy
*
FnIP	2	110	Vmeas5	0.7071068
Vmeas5	31	110	dc	0
VnIP	30	110	dc	0.65
DnIP	30	31	DIPnoisy
FnIP1	110	2	Vmeas6	0.7071068
Vmeas6	33	110	dc	0
VnIP1	32	110	dc	0.65
DnIP1	32	33	DIPnoisy
*
*
***CMRR***
RcmrrP	3	10	Rideal	1e12
RcmrrN	10	9	Rideal	1e12
g10	11	110	10	110	-1e-10
Lcmrr	11	12	1e-12
Rcmrr	12	110	Rideal	1e3
e4	5	3	11	110	1
*
*
***Power Down***
VPD	111	80	dc	1
VPD1	81	0	dc	0.2
RPD	111	106	Rideal	1e6
ePD	80	113	82	0	1
RDP1	82	0	Rideal	1e3
CPD	82	0	1e-10
S5	81	82	83	113	Switch
CDP1	83	0	1e-12
RPD2	106	83	1e6
*
*
***Gain Split***
g200	200	110	7	9	1
R200	200	110	Rideal	1e5
*
*
***Dominant Pole at 0.7 Hz***
g210	210	110	Value={limit(V(200,110)*1.39e-5,.1403,-.1403)}
R210	210	110	Rideal	2.275e6
C210	210	110	1e-7
*
*
***Output Voltage Clamp-1***
RX2	60	210	Rideal	0.001
DzVoutP	61	60	DzVoutP
DzVoutN	60	62	DzVoutN
DVoutP	61	63	diode
DVoutN	64	62	diode
VoutP	65	63	dc	6.5
VoutN	64	66	dc	5.1
e60	65	110	111	110	1.0024
e61	66	110	112	110	1.0024
*
*
***Pole at 11MHz***
g220	220	110	210	110	0.001
R220	220	110	Rideal	1000
C220	220	110	14.4686e-12
*
***Pole at 14MHz***
g230	230	110	220	110	0.001
R230	230	110	Rideal	1000
C230	230	110	11.3682e-12
*
***Buffer***
g240	240	110	230	110	0.001
R240	240	110	Rideal	1000
*
***Buffer***
g245	245	110	240	110	0.001
R245	245	110	Rideal	1000
*
***Buffer***
g250	250	110	245	110	0.001
R250	250	110	Rideal	1000
*
***Buffer***
g255	255	110	250	110	0.001
R255	255	110	Rideal	1000
*
***Buffer***
g260	260	110	255	110	0.001
R260	260	110	Rideal	1000
*
***Buffer***
g265	265	110	260	110	0.001
R265	265	110	Rideal	1000
*
***Buffer***
g270	270	110	265	110	0.001
R270	270	110	Rideal	1000
*
***Buffer***
R281	285	110	Rideal	1E6
R280	280	285	Rideal	100
e280	280	110	270	110	1
*
***Peak: f=3.5MHz, Zeta=0.7, Gain=2.4dB***
e290	290	110	285	110	1
L290	290	291	324.806e-9
C290	291	292	6366.191e-12
R291	292	110	Rideal	31.421
e295	295	110	292	110	1.3183
R290	290	292	Rideal	10
*
*
***Output Stage***
g300	300	110	295	110	0.001
R300	300	110	Rideal	1000
e301	301	110	300	110	1
Rout	302	303	Rideal	 90
Lout	303	310	3700e-9
Cout	310	110	16e-12
*
*
***Output Current Limit***
H1	301	304	Vsense1	100
Vsense1	301	302	dc	0
VIoutP	305	304	dc	0.836
VIoutN	304	306	dc	2.336
DIoutP	307	305	diode
DIoutN	306	307	diode
Rx3	307	300	Rideal	0.001
*
*
***Output Clamp-2***
VoutP1	111	73	dc	2.185
VoutN1	74	112	dc	0.785
DVoutP1	75	73	diode
DVoutN1	74	75	diode
RX4	75	310	Rideal	0.001
*
*
***Supply Currents***
FIoVcc	314	110	Vmeas8	1
Vmeas8	310	311	dc	0
R314	110	314	Rideal	1e9
DzOVcc	110	314	diode
DOVcc	102	314	diode
RX5	311	312	Rideal	0.001
FIoVee	315	110	Vmeas9	1
Vmeas9	312	313	dc	0
R315	315	110	Rideal	1e9
DzOVee	315	110	diode
DOVee	315	103	diode
*
*
***Output Switch***
S4	104	313	106	113	Switch
*
*
*** Common Models ***
.model	diode	d(bv=100)
.model	Switch	vswitch(Von=0.205,Voff=0.195,ron=10,roff=1e6)
.model	Sswitch	vswitch(Von=4.5,Voff=0.1,ron=1000,roff=1e6)
.model	DzVoutP	D(BV=4.3)
.model	DzVoutN	D(BV=4.3)
.model	DVnoisy	D(IS=7.28e-15 KF=8.83e-17)
.model	DINnoisy	D(IS=1.73e-25 KF=2.51e-21)
.model	DIPnoisy	D(IS=1.73e-25 KF=2.51e-21)
.model	Rideal	res(T_ABS=-273)
*
.ends Buffer
*
.ends ADA4530